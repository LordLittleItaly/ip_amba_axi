
`include "ip_amba_axi_top_defines.vh"
`include "ip_amba_axi_top_parameters.vh"

module ip_amba_axi_master_top `IP_AMBA_AXI_PARAM_DECL (  

    // AHB Interface Side Signals
    // Global Inputs
    
    // -------------
    // Master Inputs
    // -------------
    
    // --------------
    // Master Outputs
    // --------------
    
    // CPU / Application Layer's End's Control Signals
    // To CPU / Application Layer ( Outputs )
    
    // From CPU / Application Layer ( Inputs )

);

endmodule
