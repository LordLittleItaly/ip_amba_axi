
// ---------------
// Feature Support
// ---------------

