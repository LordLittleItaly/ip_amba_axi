// *******************************************************
// Date Created   : 18 January, 2020
// Author         : :P
// *******************************************************

// Declaration Parameters
// ----------------------
`define IP_AMBA_AXI_PARAM_DECL      #( )
